LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GUTI_ALU IS 
	PORT(STORING_CLOCK,
		  RUNNING_CLOCK,
		  STORE_SIGNAL,SAVINGEVALUATING :IN STD_LOGIC;
		REGISTER_ONE_ADDRESS,REGISTER_TWO_ADDRESS,COMPUTATION_RESULT:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	COMPLETEINSTRUCTION,RAMTEMPORARY_DATA: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_IN_REGISTER_ONE,DATA_IN_REGISTER_TWO,COMPLETERESULT:OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END GUTI_ALU;

ARCHITECTURE DESIGN OF GUTI_ALU IS

	COMPONENT GUTI_INSTRUCTION_INTERPRETATION IS 
		PORT( PERFORMANCECLOCK: IN STD_LOGIC;
		OPERATION: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		WORDONE, WORDTWO: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		COMPUTATION: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;

	COMPONENT GUTI_3_PORT_MEMORY IS
		PORT
		(	CLOCK: IN STD_LOGIC ;
			DATA: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			RDADDRESS_A: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			RDADDRESS_B: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			WRADDRESS: IN STD_LOGIC_VECTOR (4 DOWNTO 0); 
			WREN: IN STD_LOGIC := '1';
			QA: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			QB: OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
	END COMPONENT;

	SIGNAL 	TEMPORARY_DATA,FINAL_OUTPUT,
				TEMPORARY_FINAL_OUTPUT,
				TEMPORARY_A,TEMPORARY_B,
				FIRST_TEMPORARY_A,
				FIRST_TEMPORARY_B,
				EXTENDEDVALUE,
				DOT_TEMP,
				DOT_COMPLETE,
				BRANCH:STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL OPCODE,TEMPORARY_OPCODE : STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL TEMPORARY_REGISTER1,
			 TEMPORARY_REGISTER2,
			 TEMPORARY_WRITE,
			 HOLD_A,
			 HOLDB,
			 HOLDWRITE,
			 WRITE_HOLD: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL IMMEDIATE16: STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL SIGNEXTENSION,HOLD_CLOCK: STD_LOGIC;
	SIGNAL ARRAY1SIZE,ARRAY2SIZE:STD_LOGIC_VECTOR(3 DOWNTO 0);

	BEGIN
		ARRAY1SIZE<=COMPLETEINSTRUCTION(6 DOWNTO 3);
		ARRAY2SIZE<=COMPLETEINSTRUCTION(10 DOWNTO 7);
		BRANCH<=EXTENDEDVALUE;
		OPCODE <= COMPLETEINSTRUCTION(31 DOWNTO 26);
		HOLD_A <= REGISTER_ONE_ADDRESS WHEN SAVINGEVALUATING='0' ELSE TEMPORARY_REGISTER1;
		HOLDB <= REGISTER_TWO_ADDRESS WHEN SAVINGEVALUATING='0' ELSE TEMPORARY_REGISTER2;
		HOLDWRITE <= COMPUTATION_RESULT WHEN SAVINGEVALUATING='0' ELSE TEMPORARY_WRITE;
		IMMEDIATE16 <= COMPLETEINSTRUCTION(15 DOWNTO 0);
		EXTENDEDVALUE(15 DOWNTO 0) <= IMMEDIATE16;
		EXTENDEDVALUE(31 DOWNTO 16) <= (OTHERS => IMMEDIATE16(15));
		DOT_TEMP<=EXTENDEDVALUE;
		
		PROCESS(OPCODE) BEGIN
			CASE OPCODE IS
				WHEN "001100" => SIGNEXTENSION<='1';
				WHEN "001110" => BRANCH<=EXTENDEDVALUE;
				WHEN "001101" =>ARRAY1SIZE<=COMPLETEINSTRUCTION(6 DOWNTO 3);
									 ARRAY2SIZE<=COMPLETEINSTRUCTION(10 DOWNTO 7);
									 DOT_COMPLETE<=DOT_TEMP;
				WHEN OTHERS=> SIGNEXTENSION<='0';
			END CASE;
		END PROCESS;
		
		TEMPORARY_REGISTER1 <= COMPLETEINSTRUCTION(25 DOWNTO 21);
		TEMPORARY_REGISTER2 <= COMPLETEINSTRUCTION(20 DOWNTO 16);
		TEMPORARY_WRITE <= COMPLETEINSTRUCTION(15 DOWNTO 11);
		
		HOLD_CLOCK <= STORING_CLOCK;
		TEMPORARY_DATA <= RAMTEMPORARY_DATA WHEN SAVINGEVALUATING = '0' ELSE FINAL_OUTPUT;
		
		
		WRITE_HOLD<=HOLDWRITE WHEN SIGNEXTENSION='0' ELSE HOLDB;
		SAVINGTO3PORTEDMEMORY:GUTI_3_PORT_MEMORY PORT MAP(HOLD_CLOCK,
											TEMPORARY_DATA,
											HOLD_A, HOLDB, WRITE_HOLD,
											STORE_SIGNAL,
											TEMPORARY_A, TEMPORARY_B);
		
		FIRST_TEMPORARY_A <= TEMPORARY_A;
		FIRST_TEMPORARY_B <= TEMPORARY_B WHEN SIGNEXTENSION='0' ELSE EXTENDEDVALUE;
		
		TEMPORARY_OPCODE <= OPCODE WHEN SIGNEXTENSION='0' ELSE "000001";
		
		INTERPRETINGTHEINSTRUCTION : GUTI_INSTRUCTION_INTERPRETATION PORT MAP(RUNNING_CLOCK,
												TEMPORARY_OPCODE,
												FIRST_TEMPORARY_A,
												FIRST_TEMPORARY_B,
												TEMPORARY_FINAL_OUTPUT);
		FINAL_OUTPUT <= TEMPORARY_FINAL_OUTPUT;
		DATA_IN_REGISTER_ONE <= TEMPORARY_A;
		DATA_IN_REGISTER_TWO <= TEMPORARY_B;
		COMPLETERESULT <=TEMPORARY_FINAL_OUTPUT;
END DESIGN;



