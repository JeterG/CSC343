//lpm_compare CBX_SINGLE_OUTPUT_FILE="ON" LPM_REPRESENTATION="SIGNED" LPM_TYPE="LPM_COMPARE" LPM_WIDTH=6 aeb agb ageb alb aleb aneb dataa datab
//VERSION_BEGIN 16.0 cbx_mgl 2016:04:20:19:36:45:SJ cbx_stratixii 2016:04:20:18:35:29:SJ cbx_util_mgl 2016:04:20:18:35:29:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463



// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
//  Your use of Altera Corporation's design tools, logic functions 
//  and other software and tools, and its AMPP partner logic 
//  functions, and any output files from any of the foregoing 
//  (including device programming or simulation files), and any 
//  associated documentation or information are expressly subject 
//  to the terms and conditions of the Altera Program License 
//  Subscription Agreement, the Altera Quartus Prime License Agreement,
//  the Altera MegaCore Function License Agreement, or other 
//  applicable license agreement, including, without limitation, 
//  that your use is for the sole purpose of programming logic 
//  devices manufactured by Altera and sold by Altera or its 
//  authorized distributors.  Please refer to the applicable 
//  agreement for further details.



//synthesis_resources = lpm_compare 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  mgm0d
	( 
	aeb,
	agb,
	ageb,
	alb,
	aleb,
	aneb,
	dataa,
	datab) /* synthesis synthesis_clearbox=1 */;
	output   aeb;
	output   agb;
	output   ageb;
	output   alb;
	output   aleb;
	output   aneb;
	input   [5:0]  dataa;
	input   [5:0]  datab;

	wire  wire_mgl_prim1_aeb;
	wire  wire_mgl_prim1_agb;
	wire  wire_mgl_prim1_ageb;
	wire  wire_mgl_prim1_alb;
	wire  wire_mgl_prim1_aleb;
	wire  wire_mgl_prim1_aneb;

	lpm_compare   mgl_prim1
	( 
	.aeb(wire_mgl_prim1_aeb),
	.agb(wire_mgl_prim1_agb),
	.ageb(wire_mgl_prim1_ageb),
	.alb(wire_mgl_prim1_alb),
	.aleb(wire_mgl_prim1_aleb),
	.aneb(wire_mgl_prim1_aneb),
	.dataa(dataa),
	.datab(datab));
	defparam
		mgl_prim1.lpm_representation = "SIGNED",
		mgl_prim1.lpm_type = "LPM_COMPARE",
		mgl_prim1.lpm_width = 6;
	assign
		aeb = wire_mgl_prim1_aeb,
		agb = wire_mgl_prim1_agb,
		ageb = wire_mgl_prim1_ageb,
		alb = wire_mgl_prim1_alb,
		aleb = wire_mgl_prim1_aleb,
		aneb = wire_mgl_prim1_aneb;
endmodule //mgm0d
//VALID FILE
