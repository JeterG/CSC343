LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY GUTI_INSTRUCTION_INTERPRETATION IS 
PORT( PERFORMANCECLOCK: IN STD_LOGIC;
		OPERATION: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		WORDONE, WORDTWO: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		COMPUTATION: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END GUTI_INSTRUCTION_INTERPRETATION;
ARCHITECTURE ARCH OF GUTI_INSTRUCTION_INTERPRETATION IS 
	BEGIN
	PROCESS(PERFORMANCECLOCK,OPERATION)
		BEGIN
			IF(PERFORMANCECLOCK = '1') THEN
				CASE OPERATION IS 
				WHEN "000000" =>
					COMPUTATION <= WORDONE AND WORDTWO;
				WHEN "000001" =>
					COMPUTATION <= WORDONE OR WORDTWO;
				WHEN "000010" =>
					COMPUTATION <= WORDONE XOR WORDTWO;
				WHEN "000011" =>
					COMPUTATION <= NOT WORDONE;
				WHEN "000100" =>
					COMPUTATION <= TO_STDLOGICVECTOR(TO_BITVECTOR(WORDONE)SLL 1);
				WHEN "000101" =>
					COMPUTATION <= TO_STDLOGICVECTOR(TO_BITVECTOR(WORDONE)SRL 1);
				WHEN "000110" =>
					COMPUTATION <= TO_STDLOGICVECTOR(TO_BITVECTOR(WORDONE)ROL 1);
				WHEN "000111" =>
					COMPUTATION <= TO_STDLOGICVECTOR(TO_BITVECTOR(WORDONE)ROR 1);
				WHEN "001000"=> IF (WORDONE<WORDTWO) THEN COMPUTATION<=WORDONE; END IF;
								  IF (WORDONE>WORDTWO) THEN COMPUTATION<=WORDTWO; END IF;
				WHEN "001001"=> COMPUTATION<=WORDONE+WORDTWO;
				WHEN "001010"=> COMPUTATION<=WORDONE-WORDTWO;
				WHEN "001011"=> COMPUTATION<=WORDONE(15 DOWNTO 0)*WORDTWO(15 DOWNTO 0);
				WHEN OTHERS =>
				NULL;
				END CASE;
			END IF;
		END PROCESS;
END ARCH;



