LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY ALTERA_MF;
USE ALTERA_MF.ALL;
ENTITY GUTI_3_PORT_MEMORY IS
PORT
(	CLOCK: IN STD_LOGIC ;
	DATA: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	RDADDRESS_A: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	RDADDRESS_B: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	WRADDRESS: IN STD_LOGIC_VECTOR (4 DOWNTO 0); 
	WREN: IN STD_LOGIC := '1';
	QA: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	QB: OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END GUTI_3_PORT_MEMORY;
ARCHITECTURE SYN OF GUTI_3_PORT_MEMORY IS
SIGNAL SUB_WIRE0: STD_LOGIC_VECTOR (31 DOWNTO 0);
SIGNAL SUB_WIRE1: STD_LOGIC_VECTOR (31 DOWNTO 0);
COMPONENT ALT3PRAM
GENERIC (INDATA_ACLR: STRING;
			INDATA_REG: STRING;
			INTENDED_DEVICE_FAMILY: STRING;
			LPM_TYPE: STRING;
			OUTDATA_ACLR_A: STRING;
			OUTDATA_ACLR_B: STRING;
			OUTDATA_REG_A: STRING;
			OUTDATA_REG_B: STRING;
			RDADDRESS_ACLR_A: STRING;
			RDADDRESS_ACLR_B: STRING;
			RDADDRESS_REG_A: STRING;
			RDADDRESS_REG_B: STRING;
			RDCONTROL_ACLR_A: STRING;
			RDCONTROL_ACLR_B: STRING;
			RDCONTROL_REG_A: STRING;
			RDCONTROL_REG_B: STRING;
			WIDTH: NATURAL;
			WIDTHAD: NATURAL;
			WRITE_ACLR: STRING;
			WRITE_REG: STRING); 
PORT (QA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		OUTCLOCK: IN STD_LOGIC ;
		QB : OUT STD_LOGIC_VECTOR (31 DOWNTO 0); 
		WREN,INCLOCK : IN STD_LOGIC ;
		DATA: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		RDADDRESS_A : IN STD_LOGIC_VECTOR (4 DOWNTO 0); 
		WRADDRESS: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		RDADDRESS_B : IN STD_LOGIC_VECTOR (4 DOWNTO 0)
);
END COMPONENT;
BEGIN
	QA<= SUB_WIRE0(31 DOWNTO 0);
	QB<= SUB_WIRE1(31 DOWNTO 0);
	ALT3PRAM_COMPONENT : ALT3PRAM
GENERIC MAP (INDATA_ACLR => "OFF", 
				INDATA_REG=> "INCLOCK",
				INTENDED_DEVICE_FAMILY => "STRATIX II", 
				LPM_TYPE =>"ALT3PRAM",
				OUTDATA_ACLR_A => "OFF", 
				OUTDATA_ACLR_B=> "OFF", 
				OUTDATA_REG_A => "OUTCLOCK",
				OUTDATA_REG_B => "OUTCLOCK",
				RDADDRESS_ACLR_A => "OFF",
				RDADDRESS_ACLR_B => "OFF",
				RDADDRESS_REG_A => "INCLOCK",
				RDADDRESS_REG_B => "INCLOCK",
				RDCONTROL_ACLR_A => "OFF",
				RDCONTROL_ACLR_B => "OFF",
				RDCONTROL_REG_A => "UNREGISTERED",
				RDCONTROL_REG_B => "UNREGISTERED", 
				WIDTH=> 32,
				WIDTHAD => 5, 
				WRITE_ACLR =>"OFF", 
				WRITE_REG =>"INCLOCK")
PORT MAP (OUTCLOCK => CLOCK, 
			WREN=> WREN, 
			INCLOCK =>CLOCK, 
			DATA => DATA,
			RDADDRESS_A => RDADDRESS_A,
			WRADDRESS => WRADDRESS,
			RDADDRESS_B => RDADDRESS_B, 
			QA =>SUB_WIRE0,
			QB => SUB_WIRE1);
END SYN;


