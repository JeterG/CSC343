Library ieee;--JETER GUTIERREZ MAY 10, 2017
use ieee.std_logic_1164.all;--JETER GUTIERREZ MAY 10, 2017
entity GUTI_hex is--JETER GUTIERREZ MAY 10, 2017
	port(--JETER GUTIERREZ MAY 10, 2017
		bi : in std_logic_vector(3 downto 0) := X"0";--JETER GUTIERREZ MAY 10, 2017
		seg : out std_logic_vector(6 downto 0) := "0000000"--JETER GUTIERREZ MAY 10, 2017
	);--JETER GUTIERREZ MAY 10, 2017
end entity;--JETER GUTIERREZ MAY 10, 2017
architecture arch of GUTI_hex is--JETER GUTIERREZ MAY 10, 2017
begin--JETER GUTIERREZ MAY 10, 2017
	with bi select--JETER GUTIERREZ MAY 10, 2017
		seg <="1000000" when "0000", --JETER GUTIERREZ MAY 10, 2017
				"1111001" when "0001", --JETER GUTIERREZ MAY 10, 2017
				"0100100" when "0010", --JETER GUTIERREZ MAY 10, 2017
				"0110000" when "0011", --JETER GUTIERREZ MAY 10, 2017
				"0011001" when "0100", --JETER GUTIERREZ MAY 10, 2017
				"0010010" when "0101", --JETER GUTIERREZ MAY 10, 2017
				"0000010" when "0110",--JETER GUTIERREZ MAY 10, 2017
				"1111000" when "0111", --JETER GUTIERREZ MAY 10, 2017
				"0000000" when "1000", --JETER GUTIERREZ MAY 10, 2017
				"0011000" when "1001", --JETER GUTIERREZ MAY 10, 2017
				"0001000" when "1010",--JETER GUTIERREZ MAY 10, 2017
				"0000011" when "1011", --JETER GUTIERREZ MAY 10, 2017
				"1000110" when "1100", --JETER GUTIERREZ MAY 10, 2017
				"0100001" when "1101", --JETER GUTIERREZ MAY 10, 2017
				"0000110" when "1110", --JETER GUTIERREZ MAY 10, 2017
				"0001110" when "1111", --JETER GUTIERREZ MAY 10, 2017
				"1111111" when others;--JETER GUTIERREZ MAY 10, 2017
end arch;--JETER GUTIERREZ MAY 10, 2017
