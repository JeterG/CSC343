library IEEE;--JETER GUTIERREZ
use IEEE.STD_LOGIC_1164.all;--JETER GUTIERREZ
entity decode4to16 is --JETER GUTIERREZ
port(--JETER GUTIERREZ
oct : in std_logic_vector(3 downto 0);--JETER GUTIERREZ
dec : out std_logic_vector(15 downto 0));--JETER GUTIERREZ
end decode4to16;--JETER GUTIERREZ
architecture arch of decode4to16 is--JETER GUTIERREZ
begin--JETER GUTIERREZ
with oct select--JETER GUTIERREZ
dec <= "0000000000000001" when "0000",--JETER GUTIERREZ
"0000000000000010" when "0001",--JETER GUTIERREZ
"0000000000000100" when "0010",--JETER GUTIERREZ
"0000000000001000" when "0011",--JETER GUTIERREZ
"0000000000010000" when "0100",--JETER GUTIERREZ
"0000000000100000" when "0101",--JETER GUTIERREZ
"0000000001000000" when "0110",--JETER GUTIERREZ
"0000000010000000" when "0111",--JETER GUTIERREZ
"0000000100000000" when "1000",--JETER GUTIERREZ
"0000001000000000" when "1001",--JETER GUTIERREZ
"0000010000000000" when "1010",--JETER GUTIERREZ
"0000100000000000" when "1011",--JETER GUTIERREZ
"0001000000000000" when "1100",--JETER GUTIERREZ
"0010000000000000" when "1101",--JETER GUTIERREZ
"0100000000000000" when "1110",--JETER GUTIERREZ
"1000000000000000" when "1111",--JETER GUTIERREZ
"0000000000000000" when others;--JETER GUTIERREZ
end arch;--JETER GUTIERREZ